`timescale 1ns / 1ps
module down_counter;
	//Inputs
	reg  clk;
	reg  reset;
	reg  [143:0] sramConfig;
	reg  [419:0] cbconfig;
	reg  [239:0] sconfig;
	reg  [8:0]   sel;
 	wire [4:0] t01;
	wire [4:0] h01;
	wire [4:0] h02;
	wire [4:0] r01;
	wire [4:0] r02;
	wire [4:0] b01;
	wire [4:0] b02;
	wire [4:0] t02;

		
	assign t01[4:0] =	5'b000zz;
	assign t02[4:0] = 5'b0;
	assign r01[4:0] = 5'b0;
	assign b02[4:0] = 5'b0;
	assign r02[4:0] = 5'b0;
	assign b01[4:0] = 5'b0;
	assign h02[4:0] = 5'b0;
	assign h01[4:0] = 5'b000zz;
	
	
	
	initial
	begin
	sramConfig = 144'b0000000000000110_0000000000000001_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000_0000000000000000;
	cbconfig   = 420'b1100000_0000011_0000101_0001001_0010001____0000000_0000000_0000000_0000000_0000000____0000000_1000100_1001000_1010000_1100000_____1010000_0000000_0000000_0000000_0000000_____0000000_0000000_0000000_0000000_0000000____0000000_0000000_0000000_0000000_0000000___0000000_0000000_0000000_0000000_0000000____0000000_0000000_0000000_0000000_0000000____0000000_0000000_0000000_0000000_0000000____0000000_0000000_0000000_0000000_0000000____0000000_0000000_0000000_0000000_0000000____0000000_0000000_0000000_0000000_0000000;
	sconfig    = 240'b00000_00000_00000_00000_00000_10000_00000_00000_00000_00000_01000_00010___00000_00000_00000_00000_00000_00000_00000_00000_00000_00000_00000_00000____00000_00000_00000_00000_00000_00000_00000_00000_00000_00000_00000_00000_____00000_00000_00000_00000_00000_00000_00000_00000_00000_00000_00000_00000;
	sel		  = 9'b111_111_111;
	end
	// Instantiate the Unit Under Test (UUT)
	fpga_seq uut (
		.clk(clk), 
		.reset(reset), 
		.sramConfig(sramConfig), 
		.cbconfig(cbconfig),
		.sconfig(sconfig), 
		.t01(t01), 
		.t02(t02), 
		.h01(h01), 
		.h02(h02), 
		.r01(r01), 
		.r02(r02), 
		.b01(b01), 
		.b02(b02),
		.sel(sel)
	);
	always
	#50 clk=~clk;
	initial begin
		// Initialize Inputs
		clk = 0;
		reset = 1;
		#5 reset = 0;
	end    
endmodule


